`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/15/2025 10:04:55 PM
// Design Name: 
// Module Name: maindec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module maindec(
    input [6:0] op,
    output [1:0] ResultSrc,
    output MemWrite,
    output Branch, ALUSrc,
    output RegWrite, Jump,
    output [1:0] ImmSrc,
    output [1:0] ALUOp
    );
    
    reg [10:0] controls;
    assign {RegWrite, ImmSrc, ALUSrc, MemWrite, ResultSrc, Branch, ALUOp, Jump} = controls;
    
    always @ (*) begin
        case (op)
            7'b0000011 : controls = 11'b1_00_1_0_01_0_00_0;     // LW
            7'b0100011 : controls = 11'b0_01_1_1_00_0_00_0;     // SW
            7'b0110011 : controls = 11'b1_xx_0_0_00_0_10_0;     // R-type (add, sub, mul, and, or, slt)
            7'b1100011 : controls = 11'b0_10_0_0_00_1_01_0;     // beq/bne
            7'b0010011 : controls = 11'b1_00_1_0_00_0_10_0;     // I-type ALU (addi, slli)
            7'b1101111 : controls = 11'b1_11_0_0_10_0_00_1;     // jal
            7'b1100111 : controls = 11'b1_00_1_0_10_0_00_1;     // jalr
            7'b1000100 : controls = 11'b0_00_0_0_00_0_11_0;     // halt - CUSTOM
            default    : controls = 11'bx_xx_x_x_xx_x_xx_x;     // Undefined
        endcase
    end
    
endmodule
